module inverter( input A, output Z);

assign Z= !A;

endmodule
